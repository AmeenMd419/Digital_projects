`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/14/2024 12:46:54 PM
// Design Name: 
// Module Name: sub_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sub_top#(S_T0=28'D131072,S_T1=28'b0_0000000000_11101100100000110,S_T2=28'D92681,S_T3=28'D50159,
S_T4=28'D0,S_T5=-28'D50159,S_T6=-28'D92681,S_T7=-28'D121094,
S_T8=-28'D131072,S_T9=-28'D121094,S_T10=-28'D92681,S_T11=-28'D50159,
S_T12=28'D0,S_T13=28'D50159,S_T14=28'D92681,S_T15=28'D121094)
                                                            (Add,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);
                                                            
                                                            
input [7:0]X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15;
output [27:0] Add;
input clk;


wire [27:0]Y0,Y1,Y2,Y3,Y4,Y5,Y6,Y7;


Decode D0(Y0,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
S_T11,S_T12,S_T13,S_T14,S_T15,X0[0],X1[0],X2[0],X3[0],X4[0],X5[0],X6[0],
X7[0],X8[0],X9[0],X10[0],X11[0],X12[0],X13[0],X14[0],X15[0],clk);

Decode D1(Y1,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
S_T11,S_T12,S_T13,S_T14,S_T15,X0[1],X1[1],X2[1],X3[1],X4[1],X5[1],X6[1],
X7[1],X8[1],X9[1],X10[1],X11[1],X12[1],X13[1],X14[1],X15[1],clk);

Decode D2(Y2,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
S_T11,S_T12,S_T13,S_T14,S_T15,X0[2],X1[2],X2[2],X3[2],X4[2],X5[2],X6[2],
X7[2],X8[2],X9[2],X10[2],X11[2],X12[2],X13[2],X14[2],X15[2],clk);

Decode D3(Y3,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
S_T11,S_T12,S_T13,S_T14,S_T15,X0[3],X1[3],X2[3],X3[3],X4[3],X5[3],X6[3],
X7[3],X8[3],X9[3],X10[3],X11[3],X12[3],X13[3],X14[3],X15[3],clk);

Decode D4(Y4,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
S_T11,S_T12,S_T13,S_T14,S_T15,X0[4],X1[4],X2[4],X3[4],X4[4],X5[4],X6[4],
X7[4],X8[4],X9[4],X10[4],X11[4],X12[4],X13[4],X14[4],X15[4],clk);

Decode D5(Y5,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
S_T11,S_T12,S_T13,S_T14,S_T15,X0[5],X1[5],X2[5],X3[5],X4[5],X5[5],X6[5],
X7[5],X8[5],X9[5],X10[5],X11[5],X12[5],X13[5],X14[5],X15[5],clk);

Decode D6(Y6,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
S_T11,S_T12,S_T13,S_T14,S_T15,X0[6],X1[6],X2[6],X3[6],X4[6],X5[6],X6[6],
X7[6],X8[6],X9[6],X10[6],X11[6],X12[6],X13[6],X14[6],X15[6],clk);

Decode D7(Y7,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
S_T11,S_T12,S_T13,S_T14,S_T15,X0[7],X1[7],X2[7],X3[7],X4[7],X5[7],X6[7],
X7[7],X8[7],X9[7],X10[7],X11[7],X12[7],X13[7],X14[7],X15[7],clk);

top T1(Add,Y0,Y1,Y2,Y3,Y4,Y5,Y6,Y7);


//Decode D8(Y8,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
//S_T11,S_T12,S_T13,S_T14,S_T15,X0[8],X1[8],X2[8],X3[8],X4[8],X5[8],X6[8],
//X7[8],X8[8],X9[8],X10[8],X11[8],X12[8],X13[8],X14[8],X15[8],clk);

//Decode D9(Y9,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
//S_T11,S_T12,S_T13,S_T14,S_T15,X0[9],X1[9],X2[9],X3[9],X4[9],X5[9],X6[9],
//X7[9],X8[9],X9[9],X10[9],X11[9],X12[9],X13[9],X14[9],X15[9],clk);

//Decode D10(Y10,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
//S_T11,S_T12,S_T13,S_T14,S_T15,X0[10],X1[10],X2[10],X3[10],X4[10],X5[10],X6[10],
//X7[10],X8[10],X9[10],X10[10],X11[10],X12[10],X13[10],X14[10],X15[10],clk);

//Decode D11(Y11,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
//S_T11,S_T12,S_T13,S_T14,S_T15,X0[11],X1[11],X2[11],X3[11],X4[11],X5[11],X6[11],
//X7[11],X8[11],X9[11],X10[11],X11[11],X12[11],X13[11],X14[11],X15[11],clk);

//Decode D12(Y12,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
//S_T11,S_T12,S_T13,S_T14,S_T15,X0[12],X1[12],X2[12],X3[12],X4[12],X5[12],X6[12],
//X7[12],X8[12],X9[12],X10[12],X11[12],X12[12],X13[12],X14[12],X15[12],clk);

//Decode D13(Y13,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
//S_T11,S_T12,S_T13,S_T14,S_T15,X0[13],X1[13],X2[13],X3[13],X4[13],X5[13],X6[13],
//X7[13],X8[13],X9[13],X10[13],X11[13],X12[13],X13[13],X14[13],X15[13],clk);

//Decode D14(Y14,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
//S_T11,S_T12,S_T13,S_T14,S_T15,X0[14],X1[14],X2[14],X3[14],X4[14],X5[14],X6[14],
//X7[14],X8[14],X9[14],X10[14],X11[14],X12[14],X13[14],X14[14],X15[14],clk);

//Decode D15(Y15,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
//S_T11,S_T12,S_T13,S_T14,S_T15,X0[15],X1[15],X2[15],X3[15],X4[15],X5[15],X6[15],
//X7[15],X8[15],X9[15],X10[15],X11[15],X12[15],X13[15],X14[15],X15[15],clk);

//Decode D16(Y16,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
//S_T11,S_T12,S_T13,S_T14,S_T15,X0[16],X1[16],X2[16],X3[16],X4[16],X5[16],X6[16],
//X7[16],X8[16],X9[16],X10[16],X11[16],X12[16],X13[16],X14[16],X15[16],clk);

//Decode D17(Y17,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
//S_T11,S_T12,S_T13,S_T14,S_T15,X0[17],X1[17],X2[17],X3[17],X4[17],X5[17],X6[17],
//X7[17],X8[17],X9[17],X10[17],X11[17],X12[17],X13[17],X14[17],X15[17],clk);

//Decode D18(Y18,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
//S_T11,S_T12,S_T13,S_T14,S_T15,X0[18],X1[18],X2[18],X3[18],X4[18],X5[18],X6[18],
//X7[18],X8[18],X9[18],X10[18],X11[18],X12[18],X13[18],X14[18],X15[18],clk);

//Decode D19(Y19,S_T0,S_T1,S_T2,S_T3,S_T4,S_T5,S_T6,S_T7,S_T8,S_T9,S_T10,
//S_T11,S_T12,S_T13,S_T14,S_T15,X0[19],X1[19],X2[19],X3[19],X4[19],X5[19],X6[19],
//X7[19],X8[19],X9[19],X10[19],X11[19],X12[19],X13[19],X14[19],X15[19],clk);

endmodule
