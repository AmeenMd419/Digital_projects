`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/16/2024 02:33:20 PM
// Design Name: 
// Module Name: super
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module super(R0,R1,R2,R3,R4,R5,R6,R7,R8,R9,R10,R11,R12,R13,R14,R15,I0,I1,I2,I3,I4,I5,I6,I7,I8,I9,I10,I11,I12,I13,I14,I15,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);
output [27:0] R0,R1,R2,R3,R4,R5,R6,R7,R8,R9,R10,R11,R12,R13,R14,R15,
I0,I1,I2,I3,I4,I5,I6,I7,I8,I9,I10,I11,I12,I13,I14,I15;
input clk;
input [7:0]X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15;

sub_top  #(.S_T0(28'D131072),.S_T1(28'D131072),
.S_T2(28'D131072),.S_T3(28'D131072),.S_T4(28'D131072),.S_T5(28'D131072),
.S_T6(28'D131072),.S_T7(28'D131072),.S_T8(28'D131072),.S_T9(28'D131072),
.S_T10(28'D131072),.S_T11(28'D131072),.S_T12(28'D131072),.S_T13(28'D131072),.S_T14(28'D131072),.S_T15(28'D131072))
                                                             S0(R0,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);


sub_top  #(.S_T0(28'D131072),.S_T1(28'D121094),
.S_T2(28'D92681),.S_T3(28'D50159),.S_T4(28'D0),.S_T5(-28'D50159),
.S_T6(-28'D92681),.S_T7(-28'D121094),.S_T8(-28'D131072),.S_T9(-28'D121094),
.S_T10(-28'D92681),.S_T11(-28'D50159),.S_T12(28'D0),.S_T13(28'D50159),.S_T14(28'D92681),.S_T15(28'D121094))
                                                             S1(R1,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);

sub_top  #(.S_T0(28'D131072),.S_T1(28'D92681),
.S_T2(28'D0),.S_T3(-28'D92681),.S_T4(-28'D131072),.S_T5(-28'D92681),
.S_T6(28'D0),.S_T7(28'D92681),.S_T8(28'D131072),.S_T9(28'D92681),
.S_T10(28'D0),.S_T11(-28'D92681),.S_T12(-28'D131072),.S_T13(-28'D92681),.S_T14(28'D0),.S_T15(28'D92681))
                                                             S2(R2,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);

sub_top  #(.S_T0(28'D131072),.S_T1(28'D50159),
.S_T2(-28'D92681),.S_T3(-28'D121094),.S_T4(28'D0),.S_T5(28'D121094),
.S_T6(28'D92681),.S_T7(-28'D50159),.S_T8(-28'D131072),.S_T9(-28'D50159),
.S_T10(28'D92681),.S_T11(28'D121094),.S_T12(28'D0),.S_T13(-28'D121094),.S_T14(-28'D92681),.S_T15(28'D50159))
                                                             S3(R3,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);


sub_top  #(.S_T0(28'D131072),.S_T1(28'D0),
.S_T2(-28'D131072),.S_T3(28'D0),.S_T4(28'D131072),.S_T5(28'D0),
.S_T6(-28'D131072),.S_T7(28'D0),.S_T8(28'D131072),.S_T9(28'D0),
.S_T10(-28'D131072),.S_T11(28'D0),.S_T12(28'D131072),.S_T13(28'D0),.S_T14(-28'D131072),.S_T15(28'D0))
                                                             S4(R4,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);

sub_top  #(.S_T0(28'D131072),.S_T1(-28'D50159),
.S_T2(-28'D92681),.S_T3(28'D121094),.S_T4(28'D0),.S_T5(-28'D121094),
.S_T6(28'D92681),.S_T7(28'D50159),.S_T8(-28'D131072),.S_T9(28'D50159),
.S_T10(28'D92681),.S_T11(-28'D121094),.S_T12(28'D0),.S_T13(28'D121094),.S_T14(-28'D92681),.S_T15(-28'D50159))
                                                             S5(R5,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);

sub_top  #(.S_T0(28'D131072),.S_T1(-28'D92681),
.S_T2(28'D0),.S_T3(28'D92681),.S_T4(-28'D131072),.S_T5(28'D92681),
.S_T6(28'D0),.S_T7(-28'D92681),.S_T8(28'D131072),.S_T9(-28'D92681),
.S_T10(28'D0),.S_T11(28'D92681),.S_T12(-28'D131072),.S_T13(28'D92681),.S_T14(28'D0),.S_T15(-28'D92681))
                                                             S6(R6,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);

sub_top  #(.S_T0(28'D131072),.S_T1(-28'D121094),
.S_T2(28'D92681),.S_T3(-28'D50159),.S_T4(28'D0),.S_T5(28'D50159),
.S_T6(-28'D92681),.S_T7(28'D121094),.S_T8(-28'D131072),.S_T9(28'D121094),
.S_T10(-28'D92681),.S_T11(28'D50159),.S_T12(28'D0),.S_T13(-28'D50159),.S_T14(28'D92681),.S_T15(-28'D121094))
                                                             S7(R7,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);
sub_top  #(.S_T0(28'D131072),.S_T1(-28'D131072),
.S_T2(28'D131072),.S_T3(-28'D131072),.S_T4(28'D131072),.S_T5(-28'D131072),
.S_T6(28'D131072),.S_T7(-28'D131072),.S_T8(28'D131072),.S_T9(-28'D131072),
.S_T10(28'D131072),.S_T11(-28'D131072),.S_T12(28'D131072),.S_T13(-28'D131072),.S_T14(28'D131072),.S_T15(-28'D131072))
                                                             S8(R8,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);
assign R9=R7; 
assign R10 =R6;
assign R11=R5;
assign R12=R4;
assign R13 =R3;
assign R14 =R2;
assign R15 =R1;
assign I0 = 0;
sub_top  #(.S_T0(28'D0),.S_T1(-28'D50159),
.S_T2(-28'D92681),.S_T3(-28'D121094),.S_T4(-28'D131072),.S_T5(-28'D121094),
.S_T6(-28'D92681),.S_T7(-28'D50159),.S_T8(-28'D0),.S_T9(28'D50159),
.S_T10(28'D92681),.S_T11(28'D121094),.S_T12(28'D131072),.S_T13(28'D121094),.S_T14(28'D92681),.S_T15(28'D50159))
                                                             K1(I1,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);
                                                             
sub_top  #(.S_T0(28'D0),.S_T1(-28'D92681),
.S_T2(-28'D131072),.S_T3(-28'D92681),.S_T4(28'D0),.S_T5(28'D92681),
.S_T6(28'D131072),.S_T7(28'D92681),.S_T8(28'D0),.S_T9(-28'D92681),
.S_T10(-28'D131072),.S_T11(-28'D92681),.S_T12(28'D0),.S_T13(28'D92681),.S_T14(28'D131072),.S_T15(28'D92681))
                                                             K2(I2,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);         

sub_top  #(.S_T0(28'D0),.S_T1(-28'D121094),
.S_T2(-28'D92681),.S_T3(28'D50159),.S_T4(28'D131072),.S_T5(28'D50159),
.S_T6(-28'D92681),.S_T7(-28'D121094),.S_T8(28'D0),.S_T9(28'D121094),
.S_T10(28'D92681),.S_T11(-28'D50159),.S_T12(-28'D131072),.S_T13(-28'D50159),.S_T14(28'D92681),.S_T15(28'D121094))
                                                             K3(I3,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);   
sub_top  #(.S_T0(28'D0),.S_T1(-28'D131072),
.S_T2(28'D0),.S_T3(28'D131072),.S_T4(28'D0),.S_T5(-28'D131072),
.S_T6(28'D0),.S_T7(28'D131072),.S_T8(28'D0),.S_T9(-28'D131072),
.S_T10(28'D0),.S_T11(28'D131072),.S_T12(28'D0),.S_T13(-28'D131072),.S_T14(28'D0),.S_T15(28'D131072))
                                                             K4(I4,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);                                                                                                                                                                           

sub_top  #(.S_T0(28'D0),.S_T1(-28'D121094),
.S_T2(28'D92681),.S_T3(28'D50159),.S_T4(-28'D131072),.S_T5(28'D50159),
.S_T6(28'D92681),.S_T7(-28'D121094),.S_T8(28'D0),.S_T9(28'D121094),
.S_T10(-28'D92681),.S_T11(-28'D50159),.S_T12(28'D131072),.S_T13(-28'D50159),.S_T14(-28'D92681),.S_T15(28'D121094))
                                                             K5(I5,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);
                                                             
sub_top  #(.S_T0(28'D0),.S_T1(-28'D92681),
.S_T2(28'D131072),.S_T3(-28'D92681),.S_T4(28'D0),.S_T5(28'D92681),
.S_T6(-28'D131072),.S_T7(28'D92681),.S_T8(28'D0),.S_T9(-28'D92681),
.S_T10(28'D131072),.S_T11(-28'D92681),.S_T12(28'D0),.S_T13(28'D92681),.S_T14(-28'D131072),.S_T15(28'D92681))
                                                             K6(I6,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);   
 
 sub_top  #(.S_T0(28'D0),.S_T1(-28'D50159),
.S_T2(28'D92681),.S_T3(-28'D121094),.S_T4(28'D131072),.S_T5(-28'D121094),
.S_T6(28'D92681),.S_T7(-28'D50159),.S_T8(28'D0),.S_T9(28'D50159),
.S_T10(-28'D92681),.S_T11(28'D121094),.S_T12(-28'D131072),.S_T13(28'D121094),.S_T14(-28'D92681),.S_T15(28'D50159))
                                                             K7(I7,X0,X1,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11,X12,X13,X14,X15,clk);  
assign I8=0;
assign I9=-I7;
assign I10=-I6;
assign I11=-I5;
assign I12=-I4;
assign I13=-I3;
assign I14=-I2;
assign I15=-I1;
                                                          
endmodule